netcdf IAPi_0000-09-01_128x256_L30_c111201 {
dimensions:
	lat = 128 ;
	lon = 256 ;
	lev = 30 ;
	ilev = 31 ;
	chars = 1 ;
	time = UNLIMITED ; // (1 currently)
variables:
	double lat(lat) ;
		lat:long_name = "latitude" ;
		lat:units = "degrees_north" ;
	double lon(lon) ;
		lon:long_name = "longitude" ;
		lon:units = "degrees_east" ;
	double lev(lev) ;
		lev:long_name = "sigma level at midpoints" ;
		lev:units = "level" ;
		lev:positive = "down" ;
		lev:standard_name = "atmosphere_sigma_pressure_coordinate" ;
	double ilev(ilev) ;
		ilev:long_name = "sigma level at interfaces" ;
		ilev:units = "level" ;
		ilev:positive = "down" ;
		ilev:standard_name = "atmosphere_sigma_pressure_coordinate" ;
	double time(time) ;
		time:long_name = "time" ;
		time:units = "days since 0010-09-01 00:00:00" ;
		time:calendar = "noleap" ;
	double gw(lat) ;
		gw:long_name = "gauss weights" ;
	double hyai(ilev) ;
		hyai:long_name = "hybrid A coefficient at layer interfaces" ;
	double hyam(lev) ;
		hyam:long_name = "hybrid A coefficient at layer midpoints" ;
	double hybi(ilev) ;
		hybi:long_name = "hybrid B coefficient at layer interfaces" ;
	double hybm(lev) ;
		hybm:long_name = "hybrid B coefficient at layer midpoints" ;
	int ndbase ;
		ndbase:long_name = "base day" ;
	int nsbase ;
		nsbase:long_name = "seconds of base day" ;
	int nbdate ;
		nbdate:long_name = "base date (YYYYMMDD)" ;
	int nbsec ;
		nbsec:long_name = "seconds of base date" ;
	int ndcur(time) ;
		ndcur:long_name = "current day (from base day)" ;
	int nscur(time) ;
		nscur:long_name = "current seconds of current day" ;
	int date(time) ;
		date:long_name = "current date (YYYYMMDD)" ;
	int datesec(time) ;
		datesec:long_name = "current seconds of current date" ;
	int nsteph(time) ;
		nsteph:long_name = "current timestep" ;
	int mdt ;
		mdt:long_name = "timestep" ;
		mdt:units = "s" ;
	int ntrk ;
		ntrk:long_name = "spectral truncation parameter K" ;
	int ntrm ;
		ntrm:long_name = "spectral truncation parameter M" ;
	int ntrn ;
		ntrn:long_name = "spectral truncation parameter N" ;
	double CWAT(time, lat, lev, lon) ;
		CWAT:long_name = "Total Grid box averaged Condensate Amount (liquid + ice)" ;
		CWAT:units = "kg/kg" ;
	double P0 ;
		P0:long_name = "reference pressure" ;
		P0:units = "Pa" ;
	double PHIS(time, lat, lon) ;
		PHIS:long_name = "Surface geopotential" ;
		PHIS:units = "m2/s2" ;
	double PS(time, lat, lon) ;
		PS:long_name = "Surface pressure" ;
		PS:units = "Pa" ;
	double Q(time, lat, lev, lon) ;
		Q:long_name = "Specific humidity" ;
		Q:units = "kg/kg" ;
	double SNOWHICE(time, lat, lon) ;
		SNOWHICE:long_name = "Water equivalent snow depth" ;
		SNOWHICE:units = "m" ;
	double T(time, lat, lev, lon) ;
		T:long_name = "Temperature" ;
		T:units = "K" ;
	double TS(time, lat, lon) ;
		TS:long_name = "Surface temperature (radiative)" ;
		TS:units = "K" ;
	double TS1(time, lat, lon) ;
		TS1:long_name = "TS1      subsoil temperature" ;
		TS1:units = "K" ;
	double TS2(time, lat, lon) ;
		TS2:long_name = "TS2      subsoil temperature" ;
		TS2:units = "K" ;
	double TS3(time, lat, lon) ;
		TS3:long_name = "TS3      subsoil temperature" ;
		TS3:units = "K" ;
	double TS4(time, lat, lon) ;
		TS4:long_name = "TS4      subsoil temperature" ;
		TS4:units = "K" ;
	double TSICE(time, lat, lon) ;
		TSICE:long_name = "Ice temperature" ;
		TSICE:units = "K" ;
	double U(time, lat, lev, lon) ;
		U:long_name = "Zonal wind" ;
		U:units = "m/s" ;
	double V(time, lat, lev, lon) ;
		V:long_name = "Meridional wind" ;
		V:units = "m/s" ;
	char date_written(time, chars) ;
	char time_written(time, chars) ;

// global attributes:
		:history = "DEC 1 2011" ;
data:

 lat = -90, -88.5826771653543, -87.1653543307087, -85.748031496063, 
    -84.3307086614173, -82.9133858267717, -81.496062992126, 
    -80.0787401574803, -78.6614173228347, -77.244094488189, 
    -75.8267716535433, -74.4094488188976, -72.992125984252, 
    -71.5748031496063, -70.1574803149606, -68.740157480315, 
    -67.3228346456693, -65.9055118110236, -64.488188976378, 
    -63.0708661417323, -61.6535433070866, -60.2362204724409, 
    -58.8188976377953, -57.4015748031496, -55.9842519685039, 
    -54.5669291338583, -53.1496062992126, -51.7322834645669, 
    -50.3149606299213, -48.8976377952756, -47.4803149606299, 
    -46.0629921259843, -44.6456692913386, -43.2283464566929, 
    -41.8110236220472, -40.3937007874016, -38.9763779527559, 
    -37.5590551181102, -36.1417322834646, -34.7244094488189, 
    -33.3070866141732, -31.8897637795276, -30.4724409448819, 
    -29.0551181102362, -27.6377952755905, -26.2204724409449, 
    -24.8031496062992, -23.3858267716535, -21.9685039370079, 
    -20.5511811023622, -19.1338582677165, -17.7165354330709, 
    -16.2992125984252, -14.8818897637795, -13.4645669291339, 
    -12.0472440944882, -10.6299212598425, -9.21259842519684, 
    -7.79527559055119, -6.37795275590551, -4.96062992125984, 
    -3.54330708661418, -2.1259842519685, -0.70866141732283, 0.70866141732283, 
    2.1259842519685, 3.54330708661418, 4.96062992125984, 6.37795275590551, 
    7.79527559055119, 9.21259842519684, 10.6299212598425, 12.0472440944882, 
    13.4645669291339, 14.8818897637795, 16.2992125984252, 17.7165354330709, 
    19.1338582677165, 20.5511811023622, 21.9685039370079, 23.3858267716535, 
    24.8031496062992, 26.2204724409449, 27.6377952755905, 29.0551181102362, 
    30.4724409448819, 31.8897637795276, 33.3070866141732, 34.7244094488189, 
    36.1417322834646, 37.5590551181102, 38.9763779527559, 40.3937007874016, 
    41.8110236220472, 43.2283464566929, 44.6456692913386, 46.0629921259843, 
    47.4803149606299, 48.8976377952756, 50.3149606299213, 51.7322834645669, 
    53.1496062992126, 54.5669291338583, 55.9842519685039, 57.4015748031496, 
    58.8188976377953, 60.2362204724409, 61.6535433070866, 63.0708661417323, 
    64.488188976378, 65.9055118110236, 67.3228346456693, 68.740157480315, 
    70.1574803149606, 71.5748031496063, 72.992125984252, 74.4094488188976, 
    75.8267716535433, 77.244094488189, 78.6614173228346, 80.0787401574803, 
    81.496062992126, 82.9133858267716, 84.3307086614173, 85.748031496063, 
    87.1653543307087, 88.5826771653543, 90 ;

 lon = 0, 1.40625, 2.8125, 4.21875, 5.625, 7.03125, 8.4375, 9.84375, 11.25, 
    12.65625, 14.0625, 15.46875, 16.875, 18.28125, 19.6875, 21.09375, 22.5, 
    23.90625, 25.3125, 26.71875, 28.125, 29.53125, 30.9375, 32.34375, 33.75, 
    35.15625, 36.5625, 37.96875, 39.375, 40.78125, 42.1875, 43.59375, 45, 
    46.40625, 47.8125, 49.21875, 50.625, 52.03125, 53.4375, 54.84375, 56.25, 
    57.65625, 59.0625, 60.46875, 61.875, 63.28125, 64.6875, 66.09375, 67.5, 
    68.90625, 70.3125, 71.71875, 73.125, 74.53125, 75.9375, 77.34375, 78.75, 
    80.15625, 81.5625, 82.96875, 84.375, 85.78125, 87.1875, 88.59375, 90, 
    91.40625, 92.8125, 94.21875, 95.625, 97.03125, 98.4375, 99.84375, 101.25, 
    102.65625, 104.0625, 105.46875, 106.875, 108.28125, 109.6875, 111.09375, 
    112.5, 113.90625, 115.3125, 116.71875, 118.125, 119.53125, 120.9375, 
    122.34375, 123.75, 125.15625, 126.5625, 127.96875, 129.375, 130.78125, 
    132.1875, 133.59375, 135, 136.40625, 137.8125, 139.21875, 140.625, 
    142.03125, 143.4375, 144.84375, 146.25, 147.65625, 149.0625, 150.46875, 
    151.875, 153.28125, 154.6875, 156.09375, 157.5, 158.90625, 160.3125, 
    161.71875, 163.125, 164.53125, 165.9375, 167.34375, 168.75, 170.15625, 
    171.5625, 172.96875, 174.375, 175.78125, 177.1875, 178.59375, 180, 
    181.40625, 182.8125, 184.21875, 185.625, 187.03125, 188.4375, 189.84375, 
    191.25, 192.65625, 194.0625, 195.46875, 196.875, 198.28125, 199.6875, 
    201.09375, 202.5, 203.90625, 205.3125, 206.71875, 208.125, 209.53125, 
    210.9375, 212.34375, 213.75, 215.15625, 216.5625, 217.96875, 219.375, 
    220.78125, 222.1875, 223.59375, 225, 226.40625, 227.8125, 229.21875, 
    230.625, 232.03125, 233.4375, 234.84375, 236.25, 237.65625, 239.0625, 
    240.46875, 241.875, 243.28125, 244.6875, 246.09375, 247.5, 248.90625, 
    250.3125, 251.71875, 253.125, 254.53125, 255.9375, 257.34375, 258.75, 
    260.15625, 261.5625, 262.96875, 264.375, 265.78125, 267.1875, 268.59375, 
    270, 271.40625, 272.8125, 274.21875, 275.625, 277.03125, 278.4375, 
    279.84375, 281.25, 282.65625, 284.0625, 285.46875, 286.875, 288.28125, 
    289.6875, 291.09375, 292.5, 293.90625, 295.3125, 296.71875, 298.125, 
    299.53125, 300.9375, 302.34375, 303.75, 305.15625, 306.5625, 307.96875, 
    309.375, 310.78125, 312.1875, 313.59375, 315, 316.40625, 317.8125, 
    319.21875, 320.625, 322.03125, 323.4375, 324.84375, 326.25, 327.65625, 
    329.0625, 330.46875, 331.875, 333.28125, 334.6875, 336.09375, 337.5, 
    338.90625, 340.3125, 341.71875, 343.125, 344.53125, 345.9375, 347.34375, 
    348.75, 350.15625, 351.5625, 352.96875, 354.375, 355.78125, 357.1875, 
    358.59375 ;

 lev = 3.64346569404006, 7.59481964632869, 14.3566322512925, 
    24.6122200042009, 38.2682997733355, 54.5954797416925, 72.0124505460262, 
    87.8212302923203, 103.317126631737, 121.547240763903, 142.994038760662, 
    168.225079774857, 197.908086702228, 232.828618958592, 273.910816758871, 
    322.241902351379, 379.100903868675, 445.992574095726, 524.687174707651, 
    609.778694808483, 691.389430314302, 763.404481112957, 820.858368650079, 
    859.53476652503, 887.020248919725, 912.644546944648, 936.198398470879, 
    957.485479535535, 976.325407391414, 992.556095123291 ;

 ilev = 2.25523952394724, 5.03169186413288, 10.1579474285245, 
    18.5553170740604, 30.6691229343414, 45.8674766123295, 63.3234828710556, 
    80.7014182209969, 94.9410423636436, 111.69321089983, 131.401270627975, 
    154.586806893349, 181.863352656364, 213.952820748091, 251.704417169094, 
    296.117216348648, 348.366588354111, 409.83521938324, 482.149928808212, 
    567.22442060709, 652.332969009876, 730.445891618729, 796.363070607185, 
    845.353666692972, 873.715866357088, 900.324631482363, 924.964462406933, 
    947.432334534824, 967.538624536246, 985.112190246582, 1000 ;

 time = 3 ;
}
